// TCES330 Spring 2025 University of Washington Tacoma Dr. Jie Sheng
// Rodney Deacon & Mahri Yalkapova
// 06-01-2025
// Week 9, Project Folder ControlUnit
// 
/*IR is purely a group of flip-flops which will 
latch out the input signal
◦ Required input signals: Clock, ld, instruction 
from instruction memory
◦ Required output signal: instruction to the finite 
state machine
*/

module IR ( input Clk, ld,
            input [15:0] inst_in,          // instruction from instruction memory
            output logic [15:0] inst_out); //instruction to the finite state machine


   always_ff @(posedge Clk) begin
      if (ld == 1) begin
         inst_out <= inst_in;
      end else begin 
         inst_out <= inst_out;
      end
   end

endmodule

// test bench
module IR_tb;

// localparams

    // wires / logic
    logic Clk, ld;
    logic [15:0] inst_in;
    logic [15:0] inst_out;

// instantiation
   IR DUT(Clk, ld, inst_in, inst_out);

   // clock
   always begin
      Clk = 0; #10;
      Clk = 1; #10;
   end

   // testbench logic
   initial begin
      ld = 1;
      inst_in = 'd444;
      
      @(posedge Clk) #1; // wait for the values to be latched
   
      assert(inst_out == 'd444)   $display("Success!!! The output should be 444, actual: %d", inst_out);
      else $error("Expecting 444, actual: %d", inst_out);

      // disable the ld, wait for sometime, test again
      @(negedge Clk) #1;
      ld = 0;
      repeat(5) @(posedge Clk) #1;
      assert(inst_out == 'd444)   $display("Success!!! The output should be 444, actual: %d", inst_out);
      else $error("Expecting 444, actual: %d", inst_out);
      

      $stop;
   end
   // monitor
   initial begin
      $monitor($realtime, " ld = %b, inst_in = %d, inst_out = %d",ld, inst_in, inst_out);
   end

endmodule
