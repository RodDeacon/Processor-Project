/*Required input signals: Clock, D_Addr, 
D_Wr, RF_s, RF_W_Addr, RF_W_en, 
RF_Ra_Addr, RF_Rb_Addr, ALU_s0
Required output signals: ALU_inA, 
ALU_inB, ALU_out*/

module Datapath#(// params
   )
   ( // input / output 
   input Clk /*input signals: Clock, D_Addr, 
D_Wr, RF_s, RF_W_Addr, RF_W_en, 
RF_Ra_Addr, RF_Rb_Addr, ALU_s0*/
      
);
// localparam

// assignments

// combinational logic

// sequential logic

// generate block

// additional logic

endmodule

module Datapath_tb();

endmodule
